module top_module (
    input clk,
    input reset,
    output OneHertz,
    output [2:0] c_enable
);
    wire [3:0] q0, q1, q2,reset_n;
    wire carry0, carry1, carry2;

    // Enable signals
    assign c_enable[0] = 1'b1;          // first counter always enabled
    assign c_enable[1] = carry0;        // second enabled on first counter rollover
    assign c_enable[2] = carry1;        // third enabled on second counter rollover
    assign reset_n = (reset | OneHertz);
    // Instantiate first BCD counter
    bcdcount counter0 (clk,reset_n,c_enable[0],q0);
    bcdcount counter1 (clk,reset_n,c_enable[1],q1);
    bcdcount counter2 (clk,reset_n,c_enable[2],q2);

    // Detect carry from first counter
    assign carry0 = (q0 == 4'd9) & c_enable[0];
    // Detect carry from second counter
    assign carry1 = (q1 == 4'd9) & c_enable[1];
    // Detect carry from third counter
    assign carry2 = (q2 == 4'd9) & c_enable[2];

    assign OneHertz = carry2;

endmodule
//From a 1000 Hz clock, derive a 1 Hz signal, called OneHertz, that could be used to drive an Enable signal for a 
//set of hour/minute/second counters to create a digital wall clock. Since we want the clock to count once per second, 
//the OneHertz signal must be asserted for exactly one cycle each second. Build the frequency divider using modulo-10 (BCD) 
//counters and as few other gates as possible. Also output the enable signals from each of the BCD counters you use 
//(c_enable[0] for the fastest counter, c_enable[2] for the slowest).